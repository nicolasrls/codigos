library ieee;
use IEEE.std_logic_1164.all;

entity div_otmz is
    port(a,b : in std_logic;
         clk, clr: in std_logic;
         resto, rst: out std_logic;
        )
end div_otmz;

architecture pdt of div_otmz is

    



end pdt;