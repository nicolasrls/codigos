library verilog;
use verilog.vl_types.all;
entity meudisplay_vlg_vec_tst is
end meudisplay_vlg_vec_tst;
