library ieee;
use IEEE.std_logic_1164.all;

entity div_notmz is
    port(a,b : in std_logic;
         clk, clr: in std_logic;
         resto, rst: out std_logic;
        )
end div_notmz;
    
architecture pdt of div_notmz is

    



end pdt;