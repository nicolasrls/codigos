library verilog;
use verilog.vl_types.all;
entity meudisplay_vlg_check_tst is
    port(
        Sa              : in     vl_logic;
        Sb              : in     vl_logic;
        Sc              : in     vl_logic;
        Sd              : in     vl_logic;
        Se              : in     vl_logic;
        Sf              : in     vl_logic;
        Sg              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end meudisplay_vlg_check_tst;
